��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  i���    V = 5      �  i���    V = 10  X 0.5      �  ii�w    
o tambien       �  ����    <2 ) Convertira Kohms a ohms recoriendo 3 zeros  a la derecha      �  I�w�    RT = 30k      �  Iy��    RT = 10k + 10k+ 10k      �  ���    1 ) Encontrar la Corriente  I      �  �.�    
I =  V / R      �  ��4�    I = 30kohms     = 30000ohms      �  	I'    I = 15 / 3000      �  	9|G    0.0005 Amperiso (Amp)      �  	Qx_    0.5 Mili amperios (mA)      �  IY�g    RT = R1 + R2 +R3 +....      �  aA�O    V / R  X  I      �  Y!�/    Ley de ohms      �  A� ��     CIRCUTIOS RESITIVOS      �  Q�    Circutio en Serie      �  iI�W    V = 10000 X 0.0005      �  i)�7    
V = I  x R                    ��� 
 CVoltmeter��  CMeter  A3O     15.0(    �� 	 CTerminal  @(A=             .@           �  @TAi              �<            4<LT     !    ��      ��  � �� �     5.00    �  � �� �              @           �  � �� �                             � �� �    %    ��      ��  � q#     5.00(     �  0X1m              $@           �  0�1�              @            $l<�     )    ��      ��  � � � �      5.00    �  �  �              .@           �  �  �              $@            � � �     -    ��      �� 	 CResistor��  CValue  � q�     10k          ��@      �?k   �  � X� m              $@����Mb@?   �  � �� �              @����Mb@�    � l� �     3    ��      ��  CBattery1�  + �S �    15V(          .@      �? V  �  ` ha }              .@����Mb@�   �  ` �a �                ����Mb@?    T |l �     8    ��      /�1�  � &� 4    10k        ��@      �?k   �  � 8� 9             $@����Mb@�   �  � 8� 9             .@����Mb@?    � 4� <    <    ��      /�1�  � �� �    10k        ��@      �?k   �  � �� �              @����Mb@?   �  � �� �                 ����Mb@�    � �� �    @    ��      /�1�  � A� O    30k          L�@      �?k   �  � (� =             .@����Mb@?   �  � T� i              �<����Mb@�    � <� T     D    ��      5�1�  + AS O    15V(          .@      �? V  �  ` (a =             .@����Mb@�   �  ` Ta i             �<����Mb@?    T <l T     H    ��                    ���  CWire  � hAi      K�  � (A)      K�  � �� �       K�  ` �� �       K�  � �� �        K�  � �� �       K�  � �� �       K�  � �� �      K�  ` �       K�  � �1�      K�  � X1Y      K�  � 8� 9      K�  � 8� 9      K�  �  � 9       K�  �  �       K�  x 8� 9      K�  ` 8y 9      K�  x  y 9       K�  x  �       K�  � �� �       K�  � 8� Y       K�  ` 8a i       K�  ` �a �        K�  ` ha �       K�  ` �� �      K�  � h� �       K�  � � )       K�  ` a )                     �                            ! M ! " " L % % R & Q & ) V ) * * U - ^ - . . Z 3 ` 3 4 4 _ 8 a 8 9 9 b < < X = [ = @ @ S A N A D f D E E e H g H I I c E " D ! O A b P N Q P & @ % R _ g f 4 * 3 ) X ` < Y Z W . Y \ = a ] ^ [ ] - U S W V \ 8 9 O I d c e L d T M T H   6        �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 